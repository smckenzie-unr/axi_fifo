library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity AXI_FIFO is
    generic(C_AXI_ADDRESS_BUS_WIDTH:)
--  Port ( );
end AXI_FIFO;

architecture synth_logic of AXI_FIFO is

begin


end synth_logic;
